`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:56:38 06/05/2018 
// Design Name: 
// Module Name:    vga 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "Definition.h"

module vga(
	clk_25M,rst,hs,vs,red,green,blue,is_snake,is_apple,is_score,is_border,is_attention,is_meditation,is_signal,x_pos,y_pos,game_status
    );
	 
	 input clk_25M,rst;
    input game_status;                           //  ������Ϸ״̬��Ϣ������ reg �ź�
	 output reg hs,vs;							  //  �У��������ź�
	 input is_signal;
	 output reg [3:0] red,green,blue;	          //  �����ɫ�ź�
	 input is_snake,is_apple;					  //  ���������ƻ��ȷ����Ϣ
	 input is_score,is_border,is_attention,is_meditation;
	 output reg [6:0] x_pos;				      //  ���x��������Ϣ�����Ϊ 640/8 = 80
	 output reg [5:0] y_pos;				      //  ���y��������Ϣ,���Ϊ 480/8 = 60
	 reg [9:0] x_pix,y_pix;
	 reg [9:0] x,y;
	 reg [9:0] x1,y1;
	 reg [9:0] x2,y2;
	 reg [9:0] x3,y3;
	 reg [9:0] x4,y4;

//	�������źţ��������źŲ���ģ��
//	640 * 480 ������Ϊ 800 * 521
	reg [9:0] hcnt = 10'd0;		//	�����ؼ���
	reg [9:0] vcnt = 10'd0;		//	�е��м���
//	reg [9:0] x,y;					//	�������������Ϣ
	parameter [9:0] 
		hcnt_max = 10'd799,
		vcnt_max = 10'd520;
	always @(posedge clk_25M or negedge rst)
	begin
		if(!rst)
			begin
			hcnt <= 10'd0;
			vcnt <= 10'd0;
			end
		else
			if(hcnt < hcnt_max)
				hcnt <= hcnt + 1;
			else
				begin
					hcnt <= 10'd0;
					if(vcnt < vcnt_max)
						vcnt <= vcnt + 1;
					else
						vcnt <= 10'd0;
				end
	end
//	�У���ͬ���źŵĲ���
//	��ʾ��������ʾǰ�ض�������Ǹߵ�ƽ�ź�
	always @ (posedge clk_25M)
	begin
		if(hcnt > 95)
			hs <= 1'b1;
		else
			hs <= 1'b0;
	end
	always @ (posedge clk_25M)
	begin
		if(vcnt > 1)
			vs <= 1'b1;
		else 
			vs <= 1'b0;
	end
//	���ɨ���������Ϣ
//	6/23 : �޸�VGA��ʾʱ��  Active Front Sync Back
//								H:	640	  16	  96   48	800
//								V:	480	  10     2   33	525
	always @ (posedge clk_25M)
	begin
		if ((hcnt > 144) && ( hcnt < 785 ) && (vcnt > 34) && (vcnt < 515))	
			begin
				x_pos <= (hcnt - 145)>>3;
				y_pos <= (vcnt - 35)>>3;
				x_pix <= hcnt - 145;
				y_pix <= vcnt - 35;
			end
		else
			begin
				x_pos <= 0;
				y_pos <= 0;
			end						
	end
//	����������ƻ��
//	����Ϊ��ɫ
//	ƻ��Ϊ��ɫ
	always @ (posedge clk_25M or negedge rst)
	begin
		if(!rst)
			{red,green,blue} <= 12'b0000_0000_0000;
		else
         if(game_status == `Start)
			begin
			if(is_snake)											//	��ɫ��
				{red,green,blue} <= 12'b1111_0000_0000;
			else if(is_apple)										//	��ɫƻ��
				{red,green,blue} <= 12'b0000_1111_0000;
			else if(is_score)										//	��ɫ����
				{red,green,blue} <= 12'b0000_0000_1111;
			else if(is_border)									//	��ɫ�߽�
				{red,green,blue} <= 12'b1111_1111_0000;
			else if(is_attention)
				{red,green,blue} <= 12'b0000_0000_1111;
			else if(is_meditation)
				{red,green,blue} <= 12'b0000_0000_1111;
			else if(is_signal)
				{red,green,blue} <= 12'b0000_0000_1111;
			else
			begin
				{red,green,blue} <= 12'b0000_0000_0000;	
				//	  �̶���ʾ������Ϣ������
				x1 <= (x_pix - 40 + 33);
				y1 <= (y_pix - 24 + 17);
				x2 <= (x_pix - 40 + 33);
				y2 <= (y_pix - 184 + 17);
				x3 <= (x_pix - 40 + 33);
				y3 <= (y_pix - 344 + 17);
				x4 <= (x_pix - 270 + 33);
				y4 <= (y_pix - 24 + 17);
			
			if(((x1==18 && y1==2)||(x1==19 && y1==2)||(x1==51 && y1==2)||(x1==52 && y1==2)||(x1==11 && y1==3)||(x1==12 && y1==3)||(x1==17 && y1==3)||(x1==18 && y1==3)||(x1==19 && y1==3)||(x1==39 && y1==3)||(x1==40 && y1==3)||(x1==41 && y1==3)||(x1==51 && y1==3)||(x1==52 && y1==3)||(x1==53 && y1==3)||(x1==10 && y1==4)||(x1==11 && y1==4)||(x1==12 && y1==4)||(x1==18 && y1==4)||(x1==19 && y1==4)||(x1==20 && y1==4)||(x1==33 && y1==4)||(x1==34 && y1==4)||(x1==35 && y1==4)||(x1==39 && y1==4)||(x1==40 && y1==4)||(x1==41 && y1==4)||(x1==45 && y1==4)||(x1==46 && y1==4)||(x1==47 && y1==4)||(x1==51 && y1==4)||(x1==52 && y1==4)||(x1==9 && y1==5)||(x1==10 && y1==5)||(x1==11 && y1==5)||(x1==18 && y1==5)||(x1==19 && y1==5)||(x1==20 && y1==5)||(x1==34 && y1==5)||(x1==35 && y1==5)||(x1==36 && y1==5)||(x1==39 && y1==5)||(x1==40 && y1==5)||(x1==41 && y1==5)||(x1==44 && y1==5)||(x1==45 && y1==5)||(x1==46 && y1==5)||(x1==51 && y1==5)||(x1==52 && y1==5)||(x1==8 && y1==6)||(x1==9 && y1==6)||(x1==10 && y1==6)||(x1==11 && y1==6)||(x1==19 && y1==6)||(x1==20 && y1==6)||(x1==21 && y1==6)||(x1==35 && y1==6)||(x1==36 && y1==6)||(x1==39 && y1==6)||(x1==40 && y1==6)||(x1==41 && y1==6)||(x1==43 && y1==6)||(x1==44 && y1==6)||(x1==45 && y1==6)||(x1==50 && y1==6)||(x1==51 && y1==6)||(x1==52 && y1==6)||(x1==8 && y1==7)||(x1==9 && y1==7)||(x1==10 && y1==7)||(x1==20 && y1==7)||(x1==21 && y1==7)||(x1==22 && y1==7)||(x1==35 && y1==7)||(x1==36 && y1==7)||(x1==39 && y1==7)||(x1==40 && y1==7)||(x1==41 && y1==7)||(x1==43 && y1==7)||(x1==44 && y1==7)||(x1==50 && y1==7)||(x1==51 && y1==7)||(x1==52 && y1==7)||(x1==7 && y1==8)||(x1==8 && y1==8)||(x1==9 && y1==8)||(x1==20 && y1==8)||(x1==21 && y1==8)||(x1==22 && y1==8)||(x1==23 && y1==8)||(x1==39 && y1==8)||(x1==40 && y1==8)||(x1==41 && y1==8)||(x1==50 && y1==8)||(x1==51 && y1==8)||(x1==52 && y1==8)||(x1==53 && y1==8)||(x1==54 && y1==8)||(x1==55 && y1==8)||(x1==56 && y1==8)||(x1==57 && y1==8)||(x1==58 && y1==8)||(x1==59 && y1==8)||(x1==60 && y1==8)||(x1==61 && y1==8)||(x1==6 && y1==9)||(x1==7 && y1==9)||(x1==8 && y1==9)||(x1==21 && y1==9)||(x1==22 && y1==9)||(x1==23 && y1==9)||(x1==24 && y1==9)||(x1==32 && y1==9)||(x1==33 && y1==9)||(x1==34 && y1==9)||(x1==35 && y1==9)||(x1==36 && y1==9)||(x1==37 && y1==9)||(x1==38 && y1==9)||(x1==39 && y1==9)||(x1==40 && y1==9)||(x1==41 && y1==9)||(x1==42 && y1==9)||(x1==43 && y1==9)||(x1==44 && y1==9)||(x1==45 && y1==9)||(x1==46 && y1==9)||(x1==49 && y1==9)||(x1==50 && y1==9)||(x1==51 && y1==9)||(x1==52 && y1==9)||(x1==53 && y1==9)||(x1==54 && y1==9)||(x1==55 && y1==9)||(x1==56 && y1==9)||(x1==57 && y1==9)||(x1==58 && y1==9)||(x1==59 && y1==9)||(x1==60 && y1==9)||(x1==5 && y1==10)||(x1==6 && y1==10)||(x1==7 && y1==10)||(x1==22 && y1==10)||(x1==23 && y1==10)||(x1==24 && y1==10)||(x1==25 && y1==10)||(x1==32 && y1==10)||(x1==33 && y1==10)||(x1==34 && y1==10)||(x1==35 && y1==10)||(x1==36 && y1==10)||(x1==37 && y1==10)||(x1==38 && y1==10)||(x1==39 && y1==10)||(x1==40 && y1==10)||(x1==41 && y1==10)||(x1==42 && y1==10)||(x1==43 && y1==10)||(x1==44 && y1==10)||(x1==45 && y1==10)||(x1==46 && y1==10)||(x1==49 && y1==10)||(x1==50 && y1==10)||(x1==57 && y1==10)||(x1==58 && y1==10)||(x1==59 && y1==10)||(x1==4 && y1==11)||(x1==5 && y1==11)||(x1==6 && y1==11)||(x1==23 && y1==11)||(x1==24 && y1==11)||(x1==25 && y1==11)||(x1==26 && y1==11)||(x1==38 && y1==11)||(x1==39 && y1==11)||(x1==40 && y1==11)||(x1==48 && y1==11)||(x1==49 && y1==11)||(x1==50 && y1==11)||(x1==57 && y1==11)||(x1==58 && y1==11)||(x1==2 && y1==12)||(x1==3 && y1==12)||(x1==4 && y1==12)||(x1==5 && y1==12)||(x1==24 && y1==12)||(x1==25 && y1==12)||(x1==26 && y1==12)||(x1==27 && y1==12)||(x1==28 && y1==12)||(x1==36 && y1==12)||(x1==37 && y1==12)||(x1==38 && y1==12)||(x1==39 && y1==12)||(x1==40 && y1==12)||(x1==41 && y1==12)||(x1==42 && y1==12)||(x1==43 && y1==12)||(x1==47 && y1==12)||(x1==48 && y1==12)||(x1==49 && y1==12)||(x1==50 && y1==12)||(x1==51 && y1==12)||(x1==57 && y1==12)||(x1==58 && y1==12)||(x1==1 && y1==13)||(x1==2 && y1==13)||(x1==3 && y1==13)||(x1==4 && y1==13)||(x1==26 && y1==13)||(x1==27 && y1==13)||(x1==28 && y1==13)||(x1==29 && y1==13)||(x1==30 && y1==13)||(x1==35 && y1==13)||(x1==36 && y1==13)||(x1==37 && y1==13)||(x1==39 && y1==13)||(x1==40 && y1==13)||(x1==41 && y1==13)||(x1==42 && y1==13)||(x1==43 && y1==13)||(x1==44 && y1==13)||(x1==47 && y1==13)||(x1==48 && y1==13)||(x1==49 && y1==13)||(x1==50 && y1==13)||(x1==51 && y1==13)||(x1==57 && y1==13)||(x1==58 && y1==13)||(x1==1 && y1==14)||(x1==2 && y1==14)||(x1==3 && y1==14)||(x1==27 && y1==14)||(x1==28 && y1==14)||(x1==29 && y1==14)||(x1==33 && y1==14)||(x1==34 && y1==14)||(x1==35 && y1==14)||(x1==36 && y1==14)||(x1==39 && y1==14)||(x1==40 && y1==14)||(x1==43 && y1==14)||(x1==44 && y1==14)||(x1==45 && y1==14)||(x1==46 && y1==14)||(x1==47 && y1==14)||(x1==48 && y1==14)||(x1==50 && y1==14)||(x1==51 && y1==14)||(x1==56 && y1==14)||(x1==57 && y1==14)||(x1==58 && y1==14)||(x1==2 && y1==15)||(x1==5 && y1==15)||(x1==6 && y1==15)||(x1==7 && y1==15)||(x1==8 && y1==15)||(x1==9 && y1==15)||(x1==10 && y1==15)||(x1==11 && y1==15)||(x1==12 && y1==15)||(x1==13 && y1==15)||(x1==14 && y1==15)||(x1==15 && y1==15)||(x1==16 && y1==15)||(x1==17 && y1==15)||(x1==18 && y1==15)||(x1==19 && y1==15)||(x1==20 && y1==15)||(x1==21 && y1==15)||(x1==22 && y1==15)||(x1==23 && y1==15)||(x1==24 && y1==15)||(x1==32 && y1==15)||(x1==33 && y1==15)||(x1==34 && y1==15)||(x1==35 && y1==15)||(x1==39 && y1==15)||(x1==40 && y1==15)||(x1==41 && y1==15)||(x1==44 && y1==15)||(x1==45 && y1==15)||(x1==46 && y1==15)||(x1==50 && y1==15)||(x1==51 && y1==15)||(x1==56 && y1==15)||(x1==57 && y1==15)||(x1==58 && y1==15)||(x1==5 && y1==16)||(x1==6 && y1==16)||(x1==7 && y1==16)||(x1==8 && y1==16)||(x1==9 && y1==16)||(x1==10 && y1==16)||(x1==11 && y1==16)||(x1==12 && y1==16)||(x1==13 && y1==16)||(x1==14 && y1==16)||(x1==15 && y1==16)||(x1==16 && y1==16)||(x1==17 && y1==16)||(x1==18 && y1==16)||(x1==19 && y1==16)||(x1==20 && y1==16)||(x1==21 && y1==16)||(x1==22 && y1==16)||(x1==23 && y1==16)||(x1==24 && y1==16)||(x1==32 && y1==16)||(x1==33 && y1==16)||(x1==39 && y1==16)||(x1==40 && y1==16)||(x1==50 && y1==16)||(x1==51 && y1==16)||(x1==56 && y1==16)||(x1==57 && y1==16)||(x1==58 && y1==16)||(x1==10 && y1==17)||(x1==11 && y1==17)||(x1==12 && y1==17)||(x1==22 && y1==17)||(x1==23 && y1==17)||(x1==24 && y1==17)||(x1==37 && y1==17)||(x1==38 && y1==17)||(x1==39 && y1==17)||(x1==50 && y1==17)||(x1==51 && y1==17)||(x1==52 && y1==17)||(x1==56 && y1==17)||(x1==57 && y1==17)||(x1==10 && y1==18)||(x1==11 && y1==18)||(x1==12 && y1==18)||(x1==22 && y1==18)||(x1==23 && y1==18)||(x1==24 && y1==18)||(x1==36 && y1==18)||(x1==37 && y1==18)||(x1==38 && y1==18)||(x1==39 && y1==18)||(x1==51 && y1==18)||(x1==52 && y1==18)||(x1==55 && y1==18)||(x1==56 && y1==18)||(x1==57 && y1==18)||(x1==10 && y1==19)||(x1==11 && y1==19)||(x1==12 && y1==19)||(x1==22 && y1==19)||(x1==23 && y1==19)||(x1==24 && y1==19)||(x1==32 && y1==19)||(x1==33 && y1==19)||(x1==34 && y1==19)||(x1==35 && y1==19)||(x1==36 && y1==19)||(x1==37 && y1==19)||(x1==38 && y1==19)||(x1==39 && y1==19)||(x1==40 && y1==19)||(x1==41 && y1==19)||(x1==42 && y1==19)||(x1==43 && y1==19)||(x1==44 && y1==19)||(x1==45 && y1==19)||(x1==46 && y1==19)||(x1==51 && y1==19)||(x1==52 && y1==19)||(x1==53 && y1==19)||(x1==55 && y1==19)||(x1==56 && y1==19)||(x1==57 && y1==19)||(x1==10 && y1==20)||(x1==11 && y1==20)||(x1==22 && y1==20)||(x1==23 && y1==20)||(x1==24 && y1==20)||(x1==32 && y1==20)||(x1==33 && y1==20)||(x1==35 && y1==20)||(x1==36 && y1==20)||(x1==37 && y1==20)||(x1==39 && y1==20)||(x1==40 && y1==20)||(x1==41 && y1==20)||(x1==42 && y1==20)||(x1==44 && y1==20)||(x1==45 && y1==20)||(x1==51 && y1==20)||(x1==52 && y1==20)||(x1==53 && y1==20)||(x1==54 && y1==20)||(x1==55 && y1==20)||(x1==56 && y1==20)||(x1==10 && y1==21)||(x1==11 && y1==21)||(x1==22 && y1==21)||(x1==23 && y1==21)||(x1==24 && y1==21)||(x1==35 && y1==21)||(x1==36 && y1==21)||(x1==44 && y1==21)||(x1==45 && y1==21)||(x1==52 && y1==21)||(x1==53 && y1==21)||(x1==54 && y1==21)||(x1==55 && y1==21)||(x1==56 && y1==21)||(x1==9 && y1==22)||(x1==10 && y1==22)||(x1==11 && y1==22)||(x1==22 && y1==22)||(x1==23 && y1==22)||(x1==34 && y1==22)||(x1==35 && y1==22)||(x1==36 && y1==22)||(x1==43 && y1==22)||(x1==44 && y1==22)||(x1==52 && y1==22)||(x1==53 && y1==22)||(x1==54 && y1==22)||(x1==55 && y1==22)||(x1==8 && y1==23)||(x1==9 && y1==23)||(x1==10 && y1==23)||(x1==22 && y1==23)||(x1==23 && y1==23)||(x1==34 && y1==23)||(x1==35 && y1==23)||(x1==36 && y1==23)||(x1==37 && y1==23)||(x1==38 && y1==23)||(x1==42 && y1==23)||(x1==43 && y1==23)||(x1==44 && y1==23)||(x1==52 && y1==23)||(x1==53 && y1==23)||(x1==54 && y1==23)||(x1==55 && y1==23)||(x1==8 && y1==24)||(x1==9 && y1==24)||(x1==10 && y1==24)||(x1==22 && y1==24)||(x1==23 && y1==24)||(x1==36 && y1==24)||(x1==37 && y1==24)||(x1==38 && y1==24)||(x1==39 && y1==24)||(x1==40 && y1==24)||(x1==41 && y1==24)||(x1==42 && y1==24)||(x1==43 && y1==24)||(x1==51 && y1==24)||(x1==52 && y1==24)||(x1==53 && y1==24)||(x1==54 && y1==24)||(x1==55 && y1==24)||(x1==56 && y1==24)||(x1==7 && y1==25)||(x1==8 && y1==25)||(x1==9 && y1==25)||(x1==21 && y1==25)||(x1==22 && y1==25)||(x1==23 && y1==25)||(x1==38 && y1==25)||(x1==39 && y1==25)||(x1==40 && y1==25)||(x1==41 && y1==25)||(x1==42 && y1==25)||(x1==43 && y1==25)||(x1==50 && y1==25)||(x1==51 && y1==25)||(x1==52 && y1==25)||(x1==53 && y1==25)||(x1==55 && y1==25)||(x1==56 && y1==25)||(x1==57 && y1==25)||(x1==5 && y1==26)||(x1==6 && y1==26)||(x1==7 && y1==26)||(x1==8 && y1==26)||(x1==21 && y1==26)||(x1==22 && y1==26)||(x1==23 && y1==26)||(x1==37 && y1==26)||(x1==38 && y1==26)||(x1==39 && y1==26)||(x1==40 && y1==26)||(x1==41 && y1==26)||(x1==42 && y1==26)||(x1==43 && y1==26)||(x1==44 && y1==26)||(x1==45 && y1==26)||(x1==49 && y1==26)||(x1==50 && y1==26)||(x1==51 && y1==26)||(x1==52 && y1==26)||(x1==56 && y1==26)||(x1==57 && y1==26)||(x1==58 && y1==26)||(x1==59 && y1==26)||(x1==3 && y1==27)||(x1==4 && y1==27)||(x1==5 && y1==27)||(x1==6 && y1==27)||(x1==7 && y1==27)||(x1==13 && y1==27)||(x1==14 && y1==27)||(x1==15 && y1==27)||(x1==16 && y1==27)||(x1==17 && y1==27)||(x1==18 && y1==27)||(x1==19 && y1==27)||(x1==20 && y1==27)||(x1==21 && y1==27)||(x1==22 && y1==27)||(x1==35 && y1==27)||(x1==36 && y1==27)||(x1==37 && y1==27)||(x1==38 && y1==27)||(x1==39 && y1==27)||(x1==42 && y1==27)||(x1==43 && y1==27)||(x1==44 && y1==27)||(x1==45 && y1==27)||(x1==48 && y1==27)||(x1==49 && y1==27)||(x1==50 && y1==27)||(x1==51 && y1==27)||(x1==57 && y1==27)||(x1==58 && y1==27)||(x1==59 && y1==27)||(x1==60 && y1==27)||(x1==2 && y1==28)||(x1==3 && y1==28)||(x1==4 && y1==28)||(x1==5 && y1==28)||(x1==6 && y1==28)||(x1==14 && y1==28)||(x1==15 && y1==28)||(x1==16 && y1==28)||(x1==17 && y1==28)||(x1==18 && y1==28)||(x1==19 && y1==28)||(x1==20 && y1==28)||(x1==21 && y1==28)||(x1==32 && y1==28)||(x1==33 && y1==28)||(x1==34 && y1==28)||(x1==35 && y1==28)||(x1==36 && y1==28)||(x1==37 && y1==28)||(x1==44 && y1==28)||(x1==46 && y1==28)||(x1==47 && y1==28)||(x1==48 && y1==28)||(x1==49 && y1==28)||(x1==50 && y1==28)||(x1==58 && y1==28)||(x1==59 && y1==28)||(x1==60 && y1==28)||(x1==61 && y1==28)||(x1==2 && y1==29)||(x1==3 && y1==29)||(x1==4 && y1==29)||(x1==32 && y1==29)||(x1==33 && y1==29)||(x1==34 && y1==29)||(x1==35 && y1==29)||(x1==47 && y1==29)||(x1==48 && y1==29)||(x1==59 && y1==29)||(x1==60 && y1==29)) ||
				// Width: 64, Height: 32 From: /home/wanncy/����/image2verilog/score.jpg
				((x2==14 && y2==2)||(x2==15 && y2==2)||(x2==16 && y2==2)||(x2==35 && y2==2)||(x2==49 && y2==2)||(x2==50 && y2==2)||(x2==51 && y2==2)||(x2==13 && y2==3)||(x2==14 && y2==3)||(x2==15 && y2==3)||(x2==34 && y2==3)||(x2==35 && y2==3)||(x2==36 && y2==3)||(x2==49 && y2==3)||(x2==50 && y2==3)||(x2==51 && y2==3)||(x2==13 && y2==4)||(x2==14 && y2==4)||(x2==15 && y2==4)||(x2==35 && y2==4)||(x2==36 && y2==4)||(x2==37 && y2==4)||(x2==38 && y2==4)||(x2==50 && y2==4)||(x2==51 && y2==4)||(x2==52 && y2==4)||(x2==12 && y2==5)||(x2==13 && y2==5)||(x2==14 && y2==5)||(x2==15 && y2==5)||(x2==36 && y2==5)||(x2==37 && y2==5)||(x2==38 && y2==5)||(x2==39 && y2==5)||(x2==51 && y2==5)||(x2==52 && y2==5)||(x2==53 && y2==5)||(x2==3 && y2==6)||(x2==4 && y2==6)||(x2==5 && y2==6)||(x2==6 && y2==6)||(x2==7 && y2==6)||(x2==8 && y2==6)||(x2==9 && y2==6)||(x2==10 && y2==6)||(x2==11 && y2==6)||(x2==12 && y2==6)||(x2==13 && y2==6)||(x2==14 && y2==6)||(x2==15 && y2==6)||(x2==16 && y2==6)||(x2==17 && y2==6)||(x2==18 && y2==6)||(x2==19 && y2==6)||(x2==20 && y2==6)||(x2==21 && y2==6)||(x2==22 && y2==6)||(x2==23 && y2==6)||(x2==24 && y2==6)||(x2==25 && y2==6)||(x2==26 && y2==6)||(x2==27 && y2==6)||(x2==28 && y2==6)||(x2==29 && y2==6)||(x2==37 && y2==6)||(x2==38 && y2==6)||(x2==39 && y2==6)||(x2==51 && y2==6)||(x2==52 && y2==6)||(x2==3 && y2==7)||(x2==4 && y2==7)||(x2==5 && y2==7)||(x2==6 && y2==7)||(x2==7 && y2==7)||(x2==8 && y2==7)||(x2==9 && y2==7)||(x2==10 && y2==7)||(x2==11 && y2==7)||(x2==12 && y2==7)||(x2==13 && y2==7)||(x2==14 && y2==7)||(x2==15 && y2==7)||(x2==16 && y2==7)||(x2==17 && y2==7)||(x2==18 && y2==7)||(x2==19 && y2==7)||(x2==20 && y2==7)||(x2==21 && y2==7)||(x2==22 && y2==7)||(x2==23 && y2==7)||(x2==24 && y2==7)||(x2==25 && y2==7)||(x2==26 && y2==7)||(x2==27 && y2==7)||(x2==28 && y2==7)||(x2==29 && y2==7)||(x2==38 && y2==7)||(x2==39 && y2==7)||(x2==42 && y2==7)||(x2==43 && y2==7)||(x2==44 && y2==7)||(x2==45 && y2==7)||(x2==46 && y2==7)||(x2==47 && y2==7)||(x2==48 && y2==7)||(x2==49 && y2==7)||(x2==50 && y2==7)||(x2==51 && y2==7)||(x2==52 && y2==7)||(x2==53 && y2==7)||(x2==54 && y2==7)||(x2==55 && y2==7)||(x2==56 && y2==7)||(x2==57 && y2==7)||(x2==58 && y2==7)||(x2==59 && y2==7)||(x2==60 && y2==7)||(x2==61 && y2==7)||(x2==11 && y2==8)||(x2==12 && y2==8)||(x2==13 && y2==8)||(x2==42 && y2==8)||(x2==43 && y2==8)||(x2==44 && y2==8)||(x2==45 && y2==8)||(x2==46 && y2==8)||(x2==47 && y2==8)||(x2==48 && y2==8)||(x2==49 && y2==8)||(x2==50 && y2==8)||(x2==51 && y2==8)||(x2==52 && y2==8)||(x2==53 && y2==8)||(x2==54 && y2==8)||(x2==55 && y2==8)||(x2==56 && y2==8)||(x2==57 && y2==8)||(x2==58 && y2==8)||(x2==59 && y2==8)||(x2==60 && y2==8)||(x2==61 && y2==8)||(x2==11 && y2==9)||(x2==12 && y2==9)||(x2==13 && y2==9)||(x2==50 && y2==9)||(x2==51 && y2==9)||(x2==52 && y2==9)||(x2==10 && y2==10)||(x2==11 && y2==10)||(x2==12 && y2==10)||(x2==33 && y2==10)||(x2==34 && y2==10)||(x2==50 && y2==10)||(x2==51 && y2==10)||(x2==52 && y2==10)||(x2==10 && y2==11)||(x2==11 && y2==11)||(x2==12 && y2==11)||(x2==33 && y2==11)||(x2==34 && y2==11)||(x2==35 && y2==11)||(x2==36 && y2==11)||(x2==50 && y2==11)||(x2==51 && y2==11)||(x2==52 && y2==11)||(x2==2 && y2==12)||(x2==3 && y2==12)||(x2==4 && y2==12)||(x2==5 && y2==12)||(x2==6 && y2==12)||(x2==7 && y2==12)||(x2==8 && y2==12)||(x2==9 && y2==12)||(x2==10 && y2==12)||(x2==11 && y2==12)||(x2==12 && y2==12)||(x2==13 && y2==12)||(x2==14 && y2==12)||(x2==15 && y2==12)||(x2==16 && y2==12)||(x2==17 && y2==12)||(x2==18 && y2==12)||(x2==19 && y2==12)||(x2==20 && y2==12)||(x2==21 && y2==12)||(x2==22 && y2==12)||(x2==23 && y2==12)||(x2==24 && y2==12)||(x2==25 && y2==12)||(x2==26 && y2==12)||(x2==27 && y2==12)||(x2==28 && y2==12)||(x2==29 && y2==12)||(x2==30 && y2==12)||(x2==31 && y2==12)||(x2==34 && y2==12)||(x2==35 && y2==12)||(x2==36 && y2==12)||(x2==37 && y2==12)||(x2==50 && y2==12)||(x2==51 && y2==12)||(x2==52 && y2==12)||(x2==2 && y2==13)||(x2==3 && y2==13)||(x2==4 && y2==13)||(x2==5 && y2==13)||(x2==6 && y2==13)||(x2==7 && y2==13)||(x2==8 && y2==13)||(x2==9 && y2==13)||(x2==10 && y2==13)||(x2==11 && y2==13)||(x2==12 && y2==13)||(x2==13 && y2==13)||(x2==14 && y2==13)||(x2==15 && y2==13)||(x2==16 && y2==13)||(x2==17 && y2==13)||(x2==18 && y2==13)||(x2==19 && y2==13)||(x2==20 && y2==13)||(x2==21 && y2==13)||(x2==22 && y2==13)||(x2==23 && y2==13)||(x2==24 && y2==13)||(x2==25 && y2==13)||(x2==26 && y2==13)||(x2==27 && y2==13)||(x2==28 && y2==13)||(x2==29 && y2==13)||(x2==30 && y2==13)||(x2==31 && y2==13)||(x2==35 && y2==13)||(x2==36 && y2==13)||(x2==37 && y2==13)||(x2==38 && y2==13)||(x2==50 && y2==13)||(x2==51 && y2==13)||(x2==52 && y2==13)||(x2==9 && y2==14)||(x2==10 && y2==14)||(x2==11 && y2==14)||(x2==36 && y2==14)||(x2==37 && y2==14)||(x2==38 && y2==14)||(x2==50 && y2==14)||(x2==51 && y2==14)||(x2==52 && y2==14)||(x2==8 && y2==15)||(x2==9 && y2==15)||(x2==10 && y2==15)||(x2==37 && y2==15)||(x2==50 && y2==15)||(x2==51 && y2==15)||(x2==52 && y2==15)||(x2==8 && y2==16)||(x2==9 && y2==16)||(x2==10 && y2==16)||(x2==43 && y2==16)||(x2==44 && y2==16)||(x2==45 && y2==16)||(x2==46 && y2==16)||(x2==47 && y2==16)||(x2==48 && y2==16)||(x2==49 && y2==16)||(x2==50 && y2==16)||(x2==51 && y2==16)||(x2==52 && y2==16)||(x2==53 && y2==16)||(x2==54 && y2==16)||(x2==55 && y2==16)||(x2==56 && y2==16)||(x2==57 && y2==16)||(x2==58 && y2==16)||(x2==59 && y2==16)||(x2==60 && y2==16)||(x2==8 && y2==17)||(x2==9 && y2==17)||(x2==43 && y2==17)||(x2==44 && y2==17)||(x2==45 && y2==17)||(x2==46 && y2==17)||(x2==47 && y2==17)||(x2==48 && y2==17)||(x2==49 && y2==17)||(x2==50 && y2==17)||(x2==51 && y2==17)||(x2==52 && y2==17)||(x2==53 && y2==17)||(x2==54 && y2==17)||(x2==55 && y2==17)||(x2==56 && y2==17)||(x2==57 && y2==17)||(x2==58 && y2==17)||(x2==59 && y2==17)||(x2==60 && y2==17)||(x2==7 && y2==18)||(x2==8 && y2==18)||(x2==9 && y2==18)||(x2==10 && y2==18)||(x2==11 && y2==18)||(x2==12 && y2==18)||(x2==13 && y2==18)||(x2==14 && y2==18)||(x2==15 && y2==18)||(x2==16 && y2==18)||(x2==17 && y2==18)||(x2==18 && y2==18)||(x2==19 && y2==18)||(x2==20 && y2==18)||(x2==21 && y2==18)||(x2==22 && y2==18)||(x2==23 && y2==18)||(x2==24 && y2==18)||(x2==25 && y2==18)||(x2==26 && y2==18)||(x2==27 && y2==18)||(x2==43 && y2==18)||(x2==44 && y2==18)||(x2==45 && y2==18)||(x2==46 && y2==18)||(x2==47 && y2==18)||(x2==48 && y2==18)||(x2==49 && y2==18)||(x2==50 && y2==18)||(x2==51 && y2==18)||(x2==52 && y2==18)||(x2==53 && y2==18)||(x2==54 && y2==18)||(x2==55 && y2==18)||(x2==56 && y2==18)||(x2==57 && y2==18)||(x2==58 && y2==18)||(x2==59 && y2==18)||(x2==60 && y2==18)||(x2==7 && y2==19)||(x2==8 && y2==19)||(x2==9 && y2==19)||(x2==10 && y2==19)||(x2==11 && y2==19)||(x2==12 && y2==19)||(x2==13 && y2==19)||(x2==14 && y2==19)||(x2==15 && y2==19)||(x2==16 && y2==19)||(x2==17 && y2==19)||(x2==18 && y2==19)||(x2==19 && y2==19)||(x2==20 && y2==19)||(x2==21 && y2==19)||(x2==22 && y2==19)||(x2==23 && y2==19)||(x2==24 && y2==19)||(x2==25 && y2==19)||(x2==26 && y2==19)||(x2==27 && y2==19)||(x2==37 && y2==19)||(x2==38 && y2==19)||(x2==51 && y2==19)||(x2==52 && y2==19)||(x2==24 && y2==20)||(x2==25 && y2==20)||(x2==26 && y2==20)||(x2==27 && y2==20)||(x2==36 && y2==20)||(x2==37 && y2==20)||(x2==38 && y2==20)||(x2==50 && y2==20)||(x2==51 && y2==20)||(x2==52 && y2==20)||(x2==23 && y2==21)||(x2==24 && y2==21)||(x2==25 && y2==21)||(x2==26 && y2==21)||(x2==36 && y2==21)||(x2==37 && y2==21)||(x2==38 && y2==21)||(x2==50 && y2==21)||(x2==51 && y2==21)||(x2==52 && y2==21)||(x2==9 && y2==22)||(x2==22 && y2==22)||(x2==23 && y2==22)||(x2==24 && y2==22)||(x2==25 && y2==22)||(x2==36 && y2==22)||(x2==37 && y2==22)||(x2==50 && y2==22)||(x2==51 && y2==22)||(x2==52 && y2==22)||(x2==8 && y2==23)||(x2==9 && y2==23)||(x2==10 && y2==23)||(x2==11 && y2==23)||(x2==21 && y2==23)||(x2==22 && y2==23)||(x2==23 && y2==23)||(x2==35 && y2==23)||(x2==36 && y2==23)||(x2==37 && y2==23)||(x2==50 && y2==23)||(x2==51 && y2==23)||(x2==52 && y2==23)||(x2==8 && y2==24)||(x2==9 && y2==24)||(x2==10 && y2==24)||(x2==11 && y2==24)||(x2==12 && y2==24)||(x2==13 && y2==24)||(x2==19 && y2==24)||(x2==20 && y2==24)||(x2==21 && y2==24)||(x2==22 && y2==24)||(x2==35 && y2==24)||(x2==36 && y2==24)||(x2==37 && y2==24)||(x2==50 && y2==24)||(x2==51 && y2==24)||(x2==52 && y2==24)||(x2==11 && y2==25)||(x2==12 && y2==25)||(x2==13 && y2==25)||(x2==14 && y2==25)||(x2==15 && y2==25)||(x2==16 && y2==25)||(x2==18 && y2==25)||(x2==19 && y2==25)||(x2==20 && y2==25)||(x2==21 && y2==25)||(x2==35 && y2==25)||(x2==36 && y2==25)||(x2==37 && y2==25)||(x2==50 && y2==25)||(x2==51 && y2==25)||(x2==52 && y2==25)||(x2==13 && y2==26)||(x2==14 && y2==26)||(x2==15 && y2==26)||(x2==16 && y2==26)||(x2==17 && y2==26)||(x2==18 && y2==26)||(x2==19 && y2==26)||(x2==20 && y2==26)||(x2==34 && y2==26)||(x2==35 && y2==26)||(x2==36 && y2==26)||(x2==50 && y2==26)||(x2==51 && y2==26)||(x2==52 && y2==26)||(x2==15 && y2==27)||(x2==16 && y2==27)||(x2==17 && y2==27)||(x2==18 && y2==27)||(x2==19 && y2==27)||(x2==20 && y2==27)||(x2==34 && y2==27)||(x2==35 && y2==27)||(x2==36 && y2==27)||(x2==40 && y2==27)||(x2==41 && y2==27)||(x2==42 && y2==27)||(x2==43 && y2==27)||(x2==44 && y2==27)||(x2==45 && y2==27)||(x2==46 && y2==27)||(x2==47 && y2==27)||(x2==48 && y2==27)||(x2==49 && y2==27)||(x2==50 && y2==27)||(x2==51 && y2==27)||(x2==52 && y2==27)||(x2==53 && y2==27)||(x2==54 && y2==27)||(x2==55 && y2==27)||(x2==56 && y2==27)||(x2==57 && y2==27)||(x2==58 && y2==27)||(x2==59 && y2==27)||(x2==60 && y2==27)||(x2==61 && y2==27)||(x2==62 && y2==27)||(x2==17 && y2==28)||(x2==18 && y2==28)||(x2==19 && y2==28)||(x2==20 && y2==28)||(x2==21 && y2==28)||(x2==22 && y2==28)||(x2==34 && y2==28)||(x2==35 && y2==28)||(x2==36 && y2==28)||(x2==40 && y2==28)||(x2==41 && y2==28)||(x2==42 && y2==28)||(x2==43 && y2==28)||(x2==44 && y2==28)||(x2==45 && y2==28)||(x2==46 && y2==28)||(x2==47 && y2==28)||(x2==48 && y2==28)||(x2==49 && y2==28)||(x2==50 && y2==28)||(x2==51 && y2==28)||(x2==52 && y2==28)||(x2==53 && y2==28)||(x2==54 && y2==28)||(x2==55 && y2==28)||(x2==56 && y2==28)||(x2==57 && y2==28)||(x2==58 && y2==28)||(x2==59 && y2==28)||(x2==60 && y2==28)||(x2==61 && y2==28)||(x2==62 && y2==28)||(x2==19 && y2==29)||(x2==20 && y2==29)||(x2==21 && y2==29)||(x2==22 && y2==29)||(x2==23 && y2==29)||(x2==33 && y2==29)||(x2==34 && y2==29)||(x2==35 && y2==29)||(x2==21 && y2==30)||(x2==22 && y2==30)||(x2==35 && y2==30)) || 
				// Width: 64, Height: 32 From: /home/wanncy/����/image2verilog/attention.png
				((x3==38 && y3==1)||(x3==39 && y3==1)||(x3==40 && y3==1)||(x3==38 && y3==2)||(x3==39 && y3==2)||(x3==40 && y3==2)||(x3==46 && y3==2)||(x3==47 && y3==2)||(x3==48 && y3==2)||(x3==49 && y3==2)||(x3==50 && y3==2)||(x3==51 && y3==2)||(x3==52 && y3==2)||(x3==53 && y3==2)||(x3==54 && y3==2)||(x3==55 && y3==2)||(x3==56 && y3==2)||(x3==57 && y3==2)||(x3==58 && y3==2)||(x3==59 && y3==2)||(x3==60 && y3==2)||(x3==2 && y3==3)||(x3==3 && y3==3)||(x3==4 && y3==3)||(x3==5 && y3==3)||(x3==6 && y3==3)||(x3==7 && y3==3)||(x3==8 && y3==3)||(x3==9 && y3==3)||(x3==10 && y3==3)||(x3==11 && y3==3)||(x3==12 && y3==3)||(x3==13 && y3==3)||(x3==14 && y3==3)||(x3==15 && y3==3)||(x3==16 && y3==3)||(x3==17 && y3==3)||(x3==18 && y3==3)||(x3==19 && y3==3)||(x3==20 && y3==3)||(x3==21 && y3==3)||(x3==22 && y3==3)||(x3==23 && y3==3)||(x3==24 && y3==3)||(x3==25 && y3==3)||(x3==26 && y3==3)||(x3==27 && y3==3)||(x3==28 && y3==3)||(x3==29 && y3==3)||(x3==30 && y3==3)||(x3==38 && y3==3)||(x3==39 && y3==3)||(x3==40 && y3==3)||(x3==46 && y3==3)||(x3==47 && y3==3)||(x3==48 && y3==3)||(x3==49 && y3==3)||(x3==50 && y3==3)||(x3==51 && y3==3)||(x3==52 && y3==3)||(x3==53 && y3==3)||(x3==54 && y3==3)||(x3==55 && y3==3)||(x3==56 && y3==3)||(x3==57 && y3==3)||(x3==58 && y3==3)||(x3==59 && y3==3)||(x3==60 && y3==3)||(x3==2 && y3==4)||(x3==3 && y3==4)||(x3==4 && y3==4)||(x3==5 && y3==4)||(x3==6 && y3==4)||(x3==7 && y3==4)||(x3==8 && y3==4)||(x3==9 && y3==4)||(x3==10 && y3==4)||(x3==11 && y3==4)||(x3==12 && y3==4)||(x3==13 && y3==4)||(x3==14 && y3==4)||(x3==15 && y3==4)||(x3==16 && y3==4)||(x3==17 && y3==4)||(x3==18 && y3==4)||(x3==19 && y3==4)||(x3==20 && y3==4)||(x3==21 && y3==4)||(x3==22 && y3==4)||(x3==23 && y3==4)||(x3==24 && y3==4)||(x3==25 && y3==4)||(x3==26 && y3==4)||(x3==27 && y3==4)||(x3==28 && y3==4)||(x3==29 && y3==4)||(x3==30 && y3==4)||(x3==38 && y3==4)||(x3==39 && y3==4)||(x3==40 && y3==4)||(x3==46 && y3==4)||(x3==47 && y3==4)||(x3==48 && y3==4)||(x3==49 && y3==4)||(x3==50 && y3==4)||(x3==51 && y3==4)||(x3==52 && y3==4)||(x3==53 && y3==4)||(x3==54 && y3==4)||(x3==55 && y3==4)||(x3==56 && y3==4)||(x3==57 && y3==4)||(x3==58 && y3==4)||(x3==59 && y3==4)||(x3==60 && y3==4)||(x3==2 && y3==5)||(x3==3 && y3==5)||(x3==4 && y3==5)||(x3==28 && y3==5)||(x3==29 && y3==5)||(x3==30 && y3==5)||(x3==38 && y3==5)||(x3==39 && y3==5)||(x3==40 && y3==5)||(x3==46 && y3==5)||(x3==47 && y3==5)||(x3==48 && y3==5)||(x3==58 && y3==5)||(x3==59 && y3==5)||(x3==60 && y3==5)||(x3==2 && y3==6)||(x3==3 && y3==6)||(x3==4 && y3==6)||(x3==28 && y3==6)||(x3==29 && y3==6)||(x3==30 && y3==6)||(x3==33 && y3==6)||(x3==34 && y3==6)||(x3==35 && y3==6)||(x3==36 && y3==6)||(x3==37 && y3==6)||(x3==38 && y3==6)||(x3==39 && y3==6)||(x3==40 && y3==6)||(x3==41 && y3==6)||(x3==42 && y3==6)||(x3==43 && y3==6)||(x3==44 && y3==6)||(x3==46 && y3==6)||(x3==47 && y3==6)||(x3==48 && y3==6)||(x3==58 && y3==6)||(x3==59 && y3==6)||(x3==60 && y3==6)||(x3==2 && y3==7)||(x3==3 && y3==7)||(x3==4 && y3==7)||(x3==7 && y3==7)||(x3==8 && y3==7)||(x3==9 && y3==7)||(x3==10 && y3==7)||(x3==11 && y3==7)||(x3==12 && y3==7)||(x3==13 && y3==7)||(x3==14 && y3==7)||(x3==15 && y3==7)||(x3==16 && y3==7)||(x3==17 && y3==7)||(x3==18 && y3==7)||(x3==19 && y3==7)||(x3==20 && y3==7)||(x3==21 && y3==7)||(x3==22 && y3==7)||(x3==23 && y3==7)||(x3==24 && y3==7)||(x3==25 && y3==7)||(x3==28 && y3==7)||(x3==29 && y3==7)||(x3==30 && y3==7)||(x3==33 && y3==7)||(x3==34 && y3==7)||(x3==35 && y3==7)||(x3==36 && y3==7)||(x3==37 && y3==7)||(x3==38 && y3==7)||(x3==39 && y3==7)||(x3==40 && y3==7)||(x3==41 && y3==7)||(x3==42 && y3==7)||(x3==43 && y3==7)||(x3==44 && y3==7)||(x3==46 && y3==7)||(x3==47 && y3==7)||(x3==48 && y3==7)||(x3==49 && y3==7)||(x3==50 && y3==7)||(x3==51 && y3==7)||(x3==52 && y3==7)||(x3==53 && y3==7)||(x3==54 && y3==7)||(x3==55 && y3==7)||(x3==56 && y3==7)||(x3==57 && y3==7)||(x3==58 && y3==7)||(x3==59 && y3==7)||(x3==60 && y3==7)||(x3==2 && y3==8)||(x3==3 && y3==8)||(x3==4 && y3==8)||(x3==6 && y3==8)||(x3==7 && y3==8)||(x3==8 && y3==8)||(x3==9 && y3==8)||(x3==10 && y3==8)||(x3==11 && y3==8)||(x3==12 && y3==8)||(x3==13 && y3==8)||(x3==14 && y3==8)||(x3==15 && y3==8)||(x3==16 && y3==8)||(x3==17 && y3==8)||(x3==18 && y3==8)||(x3==19 && y3==8)||(x3==20 && y3==8)||(x3==21 && y3==8)||(x3==22 && y3==8)||(x3==23 && y3==8)||(x3==24 && y3==8)||(x3==25 && y3==8)||(x3==26 && y3==8)||(x3==28 && y3==8)||(x3==29 && y3==8)||(x3==30 && y3==8)||(x3==38 && y3==8)||(x3==39 && y3==8)||(x3==40 && y3==8)||(x3==46 && y3==8)||(x3==47 && y3==8)||(x3==48 && y3==8)||(x3==49 && y3==8)||(x3==50 && y3==8)||(x3==51 && y3==8)||(x3==52 && y3==8)||(x3==53 && y3==8)||(x3==54 && y3==8)||(x3==55 && y3==8)||(x3==56 && y3==8)||(x3==57 && y3==8)||(x3==58 && y3==8)||(x3==59 && y3==8)||(x3==60 && y3==8)||(x3==3 && y3==9)||(x3==6 && y3==9)||(x3==7 && y3==9)||(x3==8 && y3==9)||(x3==9 && y3==9)||(x3==10 && y3==9)||(x3==11 && y3==9)||(x3==12 && y3==9)||(x3==13 && y3==9)||(x3==14 && y3==9)||(x3==15 && y3==9)||(x3==16 && y3==9)||(x3==17 && y3==9)||(x3==18 && y3==9)||(x3==19 && y3==9)||(x3==20 && y3==9)||(x3==21 && y3==9)||(x3==22 && y3==9)||(x3==23 && y3==9)||(x3==24 && y3==9)||(x3==25 && y3==9)||(x3==26 && y3==9)||(x3==37 && y3==9)||(x3==38 && y3==9)||(x3==39 && y3==9)||(x3==40 && y3==9)||(x3==46 && y3==9)||(x3==47 && y3==9)||(x3==48 && y3==9)||(x3==58 && y3==9)||(x3==59 && y3==9)||(x3==60 && y3==9)||(x3==6 && y3==10)||(x3==7 && y3==10)||(x3==8 && y3==10)||(x3==24 && y3==10)||(x3==25 && y3==10)||(x3==26 && y3==10)||(x3==37 && y3==10)||(x3==38 && y3==10)||(x3==39 && y3==10)||(x3==40 && y3==10)||(x3==41 && y3==10)||(x3==46 && y3==10)||(x3==47 && y3==10)||(x3==48 && y3==10)||(x3==58 && y3==10)||(x3==59 && y3==10)||(x3==60 && y3==10)||(x3==6 && y3==11)||(x3==7 && y3==11)||(x3==8 && y3==11)||(x3==24 && y3==11)||(x3==25 && y3==11)||(x3==26 && y3==11)||(x3==36 && y3==11)||(x3==37 && y3==11)||(x3==38 && y3==11)||(x3==39 && y3==11)||(x3==40 && y3==11)||(x3==41 && y3==11)||(x3==42 && y3==11)||(x3==43 && y3==11)||(x3==46 && y3==11)||(x3==47 && y3==11)||(x3==48 && y3==11)||(x3==58 && y3==11)||(x3==59 && y3==11)||(x3==60 && y3==11)||(x3==6 && y3==12)||(x3==7 && y3==12)||(x3==8 && y3==12)||(x3==9 && y3==12)||(x3==10 && y3==12)||(x3==11 && y3==12)||(x3==12 && y3==12)||(x3==13 && y3==12)||(x3==14 && y3==12)||(x3==15 && y3==12)||(x3==16 && y3==12)||(x3==17 && y3==12)||(x3==18 && y3==12)||(x3==19 && y3==12)||(x3==20 && y3==12)||(x3==21 && y3==12)||(x3==22 && y3==12)||(x3==23 && y3==12)||(x3==24 && y3==12)||(x3==25 && y3==12)||(x3==26 && y3==12)||(x3==36 && y3==12)||(x3==37 && y3==12)||(x3==38 && y3==12)||(x3==39 && y3==12)||(x3==40 && y3==12)||(x3==42 && y3==12)||(x3==43 && y3==12)||(x3==44 && y3==12)||(x3==46 && y3==12)||(x3==47 && y3==12)||(x3==48 && y3==12)||(x3==49 && y3==12)||(x3==50 && y3==12)||(x3==51 && y3==12)||(x3==52 && y3==12)||(x3==53 && y3==12)||(x3==54 && y3==12)||(x3==55 && y3==12)||(x3==56 && y3==12)||(x3==57 && y3==12)||(x3==58 && y3==12)||(x3==59 && y3==12)||(x3==60 && y3==12)||(x3==6 && y3==13)||(x3==7 && y3==13)||(x3==8 && y3==13)||(x3==9 && y3==13)||(x3==10 && y3==13)||(x3==11 && y3==13)||(x3==12 && y3==13)||(x3==13 && y3==13)||(x3==14 && y3==13)||(x3==15 && y3==13)||(x3==16 && y3==13)||(x3==17 && y3==13)||(x3==18 && y3==13)||(x3==19 && y3==13)||(x3==20 && y3==13)||(x3==21 && y3==13)||(x3==22 && y3==13)||(x3==23 && y3==13)||(x3==24 && y3==13)||(x3==25 && y3==13)||(x3==26 && y3==13)||(x3==35 && y3==13)||(x3==36 && y3==13)||(x3==38 && y3==13)||(x3==39 && y3==13)||(x3==40 && y3==13)||(x3==43 && y3==13)||(x3==44 && y3==13)||(x3==46 && y3==13)||(x3==47 && y3==13)||(x3==48 && y3==13)||(x3==49 && y3==13)||(x3==50 && y3==13)||(x3==51 && y3==13)||(x3==52 && y3==13)||(x3==53 && y3==13)||(x3==54 && y3==13)||(x3==55 && y3==13)||(x3==56 && y3==13)||(x3==57 && y3==13)||(x3==58 && y3==13)||(x3==59 && y3==13)||(x3==60 && y3==13)||(x3==6 && y3==14)||(x3==7 && y3==14)||(x3==8 && y3==14)||(x3==24 && y3==14)||(x3==25 && y3==14)||(x3==26 && y3==14)||(x3==34 && y3==14)||(x3==35 && y3==14)||(x3==36 && y3==14)||(x3==38 && y3==14)||(x3==39 && y3==14)||(x3==40 && y3==14)||(x3==43 && y3==14)||(x3==46 && y3==14)||(x3==47 && y3==14)||(x3==48 && y3==14)||(x3==58 && y3==14)||(x3==59 && y3==14)||(x3==60 && y3==14)||(x3==6 && y3==15)||(x3==7 && y3==15)||(x3==8 && y3==15)||(x3==24 && y3==15)||(x3==25 && y3==15)||(x3==26 && y3==15)||(x3==33 && y3==15)||(x3==34 && y3==15)||(x3==35 && y3==15)||(x3==38 && y3==15)||(x3==39 && y3==15)||(x3==40 && y3==15)||(x3==46 && y3==15)||(x3==47 && y3==15)||(x3==48 && y3==15)||(x3==58 && y3==15)||(x3==59 && y3==15)||(x3==60 && y3==15)||(x3==6 && y3==16)||(x3==7 && y3==16)||(x3==8 && y3==16)||(x3==24 && y3==16)||(x3==25 && y3==16)||(x3==26 && y3==16)||(x3==33 && y3==16)||(x3==34 && y3==16)||(x3==35 && y3==16)||(x3==38 && y3==16)||(x3==39 && y3==16)||(x3==40 && y3==16)||(x3==46 && y3==16)||(x3==47 && y3==16)||(x3==48 && y3==16)||(x3==58 && y3==16)||(x3==59 && y3==16)||(x3==60 && y3==16)||(x3==6 && y3==17)||(x3==7 && y3==17)||(x3==8 && y3==17)||(x3==9 && y3==17)||(x3==10 && y3==17)||(x3==11 && y3==17)||(x3==12 && y3==17)||(x3==13 && y3==17)||(x3==14 && y3==17)||(x3==15 && y3==17)||(x3==16 && y3==17)||(x3==17 && y3==17)||(x3==18 && y3==17)||(x3==19 && y3==17)||(x3==20 && y3==17)||(x3==21 && y3==17)||(x3==22 && y3==17)||(x3==23 && y3==17)||(x3==24 && y3==17)||(x3==25 && y3==17)||(x3==26 && y3==17)||(x3==33 && y3==17)||(x3==34 && y3==17)||(x3==38 && y3==17)||(x3==39 && y3==17)||(x3==40 && y3==17)||(x3==46 && y3==17)||(x3==47 && y3==17)||(x3==48 && y3==17)||(x3==49 && y3==17)||(x3==50 && y3==17)||(x3==51 && y3==17)||(x3==52 && y3==17)||(x3==53 && y3==17)||(x3==54 && y3==17)||(x3==55 && y3==17)||(x3==56 && y3==17)||(x3==57 && y3==17)||(x3==58 && y3==17)||(x3==59 && y3==17)||(x3==60 && y3==17)||(x3==6 && y3==18)||(x3==7 && y3==18)||(x3==8 && y3==18)||(x3==9 && y3==18)||(x3==10 && y3==18)||(x3==11 && y3==18)||(x3==12 && y3==18)||(x3==13 && y3==18)||(x3==14 && y3==18)||(x3==15 && y3==18)||(x3==16 && y3==18)||(x3==17 && y3==18)||(x3==18 && y3==18)||(x3==19 && y3==18)||(x3==20 && y3==18)||(x3==21 && y3==18)||(x3==22 && y3==18)||(x3==23 && y3==18)||(x3==24 && y3==18)||(x3==25 && y3==18)||(x3==26 && y3==18)||(x3==38 && y3==18)||(x3==39 && y3==18)||(x3==40 && y3==18)||(x3==46 && y3==18)||(x3==47 && y3==18)||(x3==48 && y3==18)||(x3==49 && y3==18)||(x3==50 && y3==18)||(x3==51 && y3==18)||(x3==52 && y3==18)||(x3==53 && y3==18)||(x3==54 && y3==18)||(x3==55 && y3==18)||(x3==56 && y3==18)||(x3==57 && y3==18)||(x3==58 && y3==18)||(x3==59 && y3==18)||(x3==60 && y3==18)||(x3==6 && y3==19)||(x3==7 && y3==19)||(x3==8 && y3==19)||(x3==15 && y3==19)||(x3==16 && y3==19)||(x3==24 && y3==19)||(x3==25 && y3==19)||(x3==26 && y3==19)||(x3==38 && y3==19)||(x3==39 && y3==19)||(x3==40 && y3==19)||(x3==46 && y3==19)||(x3==47 && y3==19)||(x3==48 && y3==19)||(x3==58 && y3==19)||(x3==59 && y3==19)||(x3==60 && y3==19)||(x3==15 && y3==20)||(x3==16 && y3==20)||(x3==17 && y3==20)||(x3==46 && y3==20)||(x3==16 && y3==21)||(x3==17 && y3==21)||(x3==41 && y3==21)||(x3==42 && y3==21)||(x3==45 && y3==21)||(x3==46 && y3==21)||(x3==47 && y3==21)||(x3==1 && y3==22)||(x3==2 && y3==22)||(x3==3 && y3==22)||(x3==4 && y3==22)||(x3==5 && y3==22)||(x3==6 && y3==22)||(x3==7 && y3==22)||(x3==8 && y3==22)||(x3==9 && y3==22)||(x3==10 && y3==22)||(x3==11 && y3==22)||(x3==12 && y3==22)||(x3==13 && y3==22)||(x3==14 && y3==22)||(x3==15 && y3==22)||(x3==16 && y3==22)||(x3==17 && y3==22)||(x3==18 && y3==22)||(x3==19 && y3==22)||(x3==20 && y3==22)||(x3==21 && y3==22)||(x3==22 && y3==22)||(x3==23 && y3==22)||(x3==24 && y3==22)||(x3==25 && y3==22)||(x3==26 && y3==22)||(x3==27 && y3==22)||(x3==28 && y3==22)||(x3==29 && y3==22)||(x3==30 && y3==22)||(x3==31 && y3==22)||(x3==35 && y3==22)||(x3==36 && y3==22)||(x3==37 && y3==22)||(x3==41 && y3==22)||(x3==42 && y3==22)||(x3==46 && y3==22)||(x3==47 && y3==22)||(x3==48 && y3==22)||(x3==57 && y3==22)||(x3==58 && y3==22)||(x3==59 && y3==22)||(x3==1 && y3==23)||(x3==2 && y3==23)||(x3==3 && y3==23)||(x3==4 && y3==23)||(x3==5 && y3==23)||(x3==6 && y3==23)||(x3==7 && y3==23)||(x3==8 && y3==23)||(x3==9 && y3==23)||(x3==10 && y3==23)||(x3==11 && y3==23)||(x3==12 && y3==23)||(x3==13 && y3==23)||(x3==14 && y3==23)||(x3==15 && y3==23)||(x3==16 && y3==23)||(x3==17 && y3==23)||(x3==18 && y3==23)||(x3==19 && y3==23)||(x3==20 && y3==23)||(x3==21 && y3==23)||(x3==22 && y3==23)||(x3==23 && y3==23)||(x3==24 && y3==23)||(x3==25 && y3==23)||(x3==26 && y3==23)||(x3==27 && y3==23)||(x3==28 && y3==23)||(x3==29 && y3==23)||(x3==30 && y3==23)||(x3==31 && y3==23)||(x3==35 && y3==23)||(x3==36 && y3==23)||(x3==37 && y3==23)||(x3==41 && y3==23)||(x3==42 && y3==23)||(x3==47 && y3==23)||(x3==48 && y3==23)||(x3==49 && y3==23)||(x3==50 && y3==23)||(x3==54 && y3==23)||(x3==58 && y3==23)||(x3==59 && y3==23)||(x3==60 && y3==23)||(x3==35 && y3==24)||(x3==36 && y3==24)||(x3==41 && y3==24)||(x3==42 && y3==24)||(x3==48 && y3==24)||(x3==49 && y3==24)||(x3==54 && y3==24)||(x3==55 && y3==24)||(x3==59 && y3==24)||(x3==60 && y3==24)||(x3==61 && y3==24)||(x3==11 && y3==25)||(x3==12 && y3==25)||(x3==20 && y3==25)||(x3==21 && y3==25)||(x3==34 && y3==25)||(x3==35 && y3==25)||(x3==36 && y3==25)||(x3==41 && y3==25)||(x3==42 && y3==25)||(x3==54 && y3==25)||(x3==55 && y3==25)||(x3==59 && y3==25)||(x3==60 && y3==25)||(x3==61 && y3==25)||(x3==9 && y3==26)||(x3==10 && y3==26)||(x3==11 && y3==26)||(x3==12 && y3==26)||(x3==19 && y3==26)||(x3==20 && y3==26)||(x3==21 && y3==26)||(x3==22 && y3==26)||(x3==23 && y3==26)||(x3==24 && y3==26)||(x3==34 && y3==26)||(x3==35 && y3==26)||(x3==41 && y3==26)||(x3==42 && y3==26)||(x3==53 && y3==26)||(x3==54 && y3==26)||(x3==55 && y3==26)||(x3==60 && y3==26)||(x3==61 && y3==26)||(x3==62 && y3==26)||(x3==6 && y3==27)||(x3==7 && y3==27)||(x3==8 && y3==27)||(x3==9 && y3==27)||(x3==10 && y3==27)||(x3==11 && y3==27)||(x3==12 && y3==27)||(x3==20 && y3==27)||(x3==21 && y3==27)||(x3==22 && y3==27)||(x3==23 && y3==27)||(x3==24 && y3==27)||(x3==25 && y3==27)||(x3==26 && y3==27)||(x3==27 && y3==27)||(x3==33 && y3==27)||(x3==34 && y3==27)||(x3==35 && y3==27)||(x3==41 && y3==27)||(x3==42 && y3==27)||(x3==53 && y3==27)||(x3==54 && y3==27)||(x3==55 && y3==27)||(x3==61 && y3==27)||(x3==3 && y3==28)||(x3==4 && y3==28)||(x3==5 && y3==28)||(x3==6 && y3==28)||(x3==7 && y3==28)||(x3==8 && y3==28)||(x3==9 && y3==28)||(x3==23 && y3==28)||(x3==24 && y3==28)||(x3==25 && y3==28)||(x3==26 && y3==28)||(x3==27 && y3==28)||(x3==28 && y3==28)||(x3==29 && y3==28)||(x3==30 && y3==28)||(x3==33 && y3==28)||(x3==34 && y3==28)||(x3==41 && y3==28)||(x3==42 && y3==28)||(x3==43 && y3==28)||(x3==44 && y3==28)||(x3==45 && y3==28)||(x3==46 && y3==28)||(x3==47 && y3==28)||(x3==48 && y3==28)||(x3==49 && y3==28)||(x3==50 && y3==28)||(x3==51 && y3==28)||(x3==52 && y3==28)||(x3==53 && y3==28)||(x3==54 && y3==28)||(x3==2 && y3==29)||(x3==3 && y3==29)||(x3==4 && y3==29)||(x3==5 && y3==29)||(x3==6 && y3==29)||(x3==7 && y3==29)||(x3==25 && y3==29)||(x3==26 && y3==29)||(x3==27 && y3==29)||(x3==28 && y3==29)||(x3==29 && y3==29)||(x3==30 && y3==29)||(x3==42 && y3==29)||(x3==43 && y3==29)||(x3==44 && y3==29)||(x3==45 && y3==29)||(x3==46 && y3==29)||(x3==47 && y3==29)||(x3==48 && y3==29)||(x3==49 && y3==29)||(x3==50 && y3==29)||(x3==51 && y3==29)||(x3==52 && y3==29)||(x3==53 && y3==29)||(x3==54 && y3==29)||(x3==2 && y3==30)||(x3==3 && y3==30)||(x3==4 && y3==30)||(x3==28 && y3==30)||(x3==29 && y3==30)||(x3==44 && y3==30)||(x3==45 && y3==30)||(x3==46 && y3==30)||(x3==47 && y3==30)||(x3==48 && y3==30)||(x3==49 && y3==30)||(x3==50 && y3==30)||(x3==51 && y3==30)) ||
				// Width: 64, Height: 32 From: /home/wanncy/����/image2verilog/dream.png
				((x4==8 && y4==1)||(x4==20 && y4==1)||(x4==8 && y4==2)||(x4==9 && y4==2)||(x4==10 && y4==2)||(x4==19 && y4==2)||(x4==20 && y4==2)||(x4==8 && y4==3)||(x4==9 && y4==3)||(x4==19 && y4==3)||(x4==20 && y4==3)||(x4==21 && y4==3)||(x4==38 && y4==3)||(x4==39 && y4==3)||(x4==40 && y4==3)||(x4==41 && y4==3)||(x4==42 && y4==3)||(x4==43 && y4==3)||(x4==44 && y4==3)||(x4==45 && y4==3)||(x4==46 && y4==3)||(x4==47 && y4==3)||(x4==48 && y4==3)||(x4==49 && y4==3)||(x4==50 && y4==3)||(x4==51 && y4==3)||(x4==52 && y4==3)||(x4==53 && y4==3)||(x4==54 && y4==3)||(x4==55 && y4==3)||(x4==56 && y4==3)||(x4==57 && y4==3)||(x4==7 && y4==4)||(x4==8 && y4==4)||(x4==9 && y4==4)||(x4==20 && y4==4)||(x4==21 && y4==4)||(x4==38 && y4==4)||(x4==39 && y4==4)||(x4==40 && y4==4)||(x4==41 && y4==4)||(x4==42 && y4==4)||(x4==43 && y4==4)||(x4==44 && y4==4)||(x4==45 && y4==4)||(x4==46 && y4==4)||(x4==47 && y4==4)||(x4==48 && y4==4)||(x4==49 && y4==4)||(x4==50 && y4==4)||(x4==51 && y4==4)||(x4==52 && y4==4)||(x4==53 && y4==4)||(x4==54 && y4==4)||(x4==55 && y4==4)||(x4==56 && y4==4)||(x4==57 && y4==4)||(x4==7 && y4==5)||(x4==8 && y4==5)||(x4==11 && y4==5)||(x4==12 && y4==5)||(x4==13 && y4==5)||(x4==14 && y4==5)||(x4==15 && y4==5)||(x4==16 && y4==5)||(x4==17 && y4==5)||(x4==18 && y4==5)||(x4==19 && y4==5)||(x4==20 && y4==5)||(x4==21 && y4==5)||(x4==22 && y4==5)||(x4==23 && y4==5)||(x4==24 && y4==5)||(x4==25 && y4==5)||(x4==26 && y4==5)||(x4==27 && y4==5)||(x4==28 && y4==5)||(x4==29 && y4==5)||(x4==30 && y4==5)||(x4==31 && y4==5)||(x4==38 && y4==5)||(x4==39 && y4==5)||(x4==56 && y4==5)||(x4==57 && y4==5)||(x4==6 && y4==6)||(x4==7 && y4==6)||(x4==8 && y4==6)||(x4==10 && y4==6)||(x4==11 && y4==6)||(x4==12 && y4==6)||(x4==13 && y4==6)||(x4==14 && y4==6)||(x4==15 && y4==6)||(x4==16 && y4==6)||(x4==17 && y4==6)||(x4==18 && y4==6)||(x4==19 && y4==6)||(x4==20 && y4==6)||(x4==21 && y4==6)||(x4==22 && y4==6)||(x4==23 && y4==6)||(x4==24 && y4==6)||(x4==25 && y4==6)||(x4==26 && y4==6)||(x4==27 && y4==6)||(x4==28 && y4==6)||(x4==29 && y4==6)||(x4==30 && y4==6)||(x4==31 && y4==6)||(x4==38 && y4==6)||(x4==39 && y4==6)||(x4==56 && y4==6)||(x4==57 && y4==6)||(x4==6 && y4==7)||(x4==7 && y4==7)||(x4==8 && y4==7)||(x4==11 && y4==7)||(x4==12 && y4==7)||(x4==13 && y4==7)||(x4==14 && y4==7)||(x4==15 && y4==7)||(x4==16 && y4==7)||(x4==17 && y4==7)||(x4==18 && y4==7)||(x4==19 && y4==7)||(x4==20 && y4==7)||(x4==21 && y4==7)||(x4==22 && y4==7)||(x4==23 && y4==7)||(x4==24 && y4==7)||(x4==25 && y4==7)||(x4==26 && y4==7)||(x4==27 && y4==7)||(x4==28 && y4==7)||(x4==29 && y4==7)||(x4==30 && y4==7)||(x4==31 && y4==7)||(x4==38 && y4==7)||(x4==39 && y4==7)||(x4==56 && y4==7)||(x4==57 && y4==7)||(x4==6 && y4==8)||(x4==7 && y4==8)||(x4==38 && y4==8)||(x4==39 && y4==8)||(x4==56 && y4==8)||(x4==57 && y4==8)||(x4==5 && y4==9)||(x4==6 && y4==9)||(x4==7 && y4==9)||(x4==38 && y4==9)||(x4==39 && y4==9)||(x4==40 && y4==9)||(x4==41 && y4==9)||(x4==42 && y4==9)||(x4==43 && y4==9)||(x4==44 && y4==9)||(x4==45 && y4==9)||(x4==46 && y4==9)||(x4==47 && y4==9)||(x4==48 && y4==9)||(x4==49 && y4==9)||(x4==50 && y4==9)||(x4==51 && y4==9)||(x4==52 && y4==9)||(x4==53 && y4==9)||(x4==54 && y4==9)||(x4==55 && y4==9)||(x4==56 && y4==9)||(x4==57 && y4==9)||(x4==5 && y4==10)||(x4==6 && y4==10)||(x4==7 && y4==10)||(x4==12 && y4==10)||(x4==13 && y4==10)||(x4==14 && y4==10)||(x4==15 && y4==10)||(x4==16 && y4==10)||(x4==17 && y4==10)||(x4==18 && y4==10)||(x4==19 && y4==10)||(x4==20 && y4==10)||(x4==21 && y4==10)||(x4==22 && y4==10)||(x4==23 && y4==10)||(x4==24 && y4==10)||(x4==25 && y4==10)||(x4==26 && y4==10)||(x4==27 && y4==10)||(x4==28 && y4==10)||(x4==29 && y4==10)||(x4==38 && y4==10)||(x4==39 && y4==10)||(x4==40 && y4==10)||(x4==41 && y4==10)||(x4==42 && y4==10)||(x4==43 && y4==10)||(x4==44 && y4==10)||(x4==45 && y4==10)||(x4==46 && y4==10)||(x4==47 && y4==10)||(x4==48 && y4==10)||(x4==49 && y4==10)||(x4==50 && y4==10)||(x4==51 && y4==10)||(x4==52 && y4==10)||(x4==53 && y4==10)||(x4==54 && y4==10)||(x4==55 && y4==10)||(x4==56 && y4==10)||(x4==57 && y4==10)||(x4==4 && y4==11)||(x4==5 && y4==11)||(x4==6 && y4==11)||(x4==7 && y4==11)||(x4==12 && y4==11)||(x4==13 && y4==11)||(x4==14 && y4==11)||(x4==15 && y4==11)||(x4==16 && y4==11)||(x4==17 && y4==11)||(x4==18 && y4==11)||(x4==19 && y4==11)||(x4==20 && y4==11)||(x4==21 && y4==11)||(x4==22 && y4==11)||(x4==23 && y4==11)||(x4==24 && y4==11)||(x4==25 && y4==11)||(x4==26 && y4==11)||(x4==27 && y4==11)||(x4==28 && y4==11)||(x4==29 && y4==11)||(x4==38 && y4==11)||(x4==39 && y4==11)||(x4==40 && y4==11)||(x4==55 && y4==11)||(x4==56 && y4==11)||(x4==57 && y4==11)||(x4==4 && y4==12)||(x4==5 && y4==12)||(x4==6 && y4==12)||(x4==7 && y4==12)||(x4==29 && y4==12)||(x4==38 && y4==12)||(x4==39 && y4==12)||(x4==56 && y4==12)||(x4==57 && y4==12)||(x4==3 && y4==13)||(x4==4 && y4==13)||(x4==5 && y4==13)||(x4==6 && y4==13)||(x4==7 && y4==13)||(x4==2 && y4==14)||(x4==3 && y4==14)||(x4==4 && y4==14)||(x4==5 && y4==14)||(x4==6 && y4==14)||(x4==7 && y4==14)||(x4==33 && y4==14)||(x4==34 && y4==14)||(x4==35 && y4==14)||(x4==36 && y4==14)||(x4==37 && y4==14)||(x4==38 && y4==14)||(x4==39 && y4==14)||(x4==40 && y4==14)||(x4==41 && y4==14)||(x4==42 && y4==14)||(x4==43 && y4==14)||(x4==44 && y4==14)||(x4==45 && y4==14)||(x4==46 && y4==14)||(x4==47 && y4==14)||(x4==48 && y4==14)||(x4==49 && y4==14)||(x4==50 && y4==14)||(x4==51 && y4==14)||(x4==52 && y4==14)||(x4==53 && y4==14)||(x4==54 && y4==14)||(x4==55 && y4==14)||(x4==56 && y4==14)||(x4==57 && y4==14)||(x4==58 && y4==14)||(x4==59 && y4==14)||(x4==60 && y4==14)||(x4==61 && y4==14)||(x4==62 && y4==14)||(x4==2 && y4==15)||(x4==3 && y4==15)||(x4==4 && y4==15)||(x4==6 && y4==15)||(x4==7 && y4==15)||(x4==12 && y4==15)||(x4==13 && y4==15)||(x4==14 && y4==15)||(x4==15 && y4==15)||(x4==16 && y4==15)||(x4==17 && y4==15)||(x4==18 && y4==15)||(x4==19 && y4==15)||(x4==20 && y4==15)||(x4==21 && y4==15)||(x4==22 && y4==15)||(x4==23 && y4==15)||(x4==24 && y4==15)||(x4==25 && y4==15)||(x4==26 && y4==15)||(x4==27 && y4==15)||(x4==28 && y4==15)||(x4==29 && y4==15)||(x4==33 && y4==15)||(x4==34 && y4==15)||(x4==35 && y4==15)||(x4==36 && y4==15)||(x4==37 && y4==15)||(x4==38 && y4==15)||(x4==39 && y4==15)||(x4==40 && y4==15)||(x4==41 && y4==15)||(x4==42 && y4==15)||(x4==43 && y4==15)||(x4==44 && y4==15)||(x4==45 && y4==15)||(x4==46 && y4==15)||(x4==47 && y4==15)||(x4==48 && y4==15)||(x4==49 && y4==15)||(x4==50 && y4==15)||(x4==51 && y4==15)||(x4==52 && y4==15)||(x4==53 && y4==15)||(x4==54 && y4==15)||(x4==55 && y4==15)||(x4==56 && y4==15)||(x4==57 && y4==15)||(x4==58 && y4==15)||(x4==59 && y4==15)||(x4==60 && y4==15)||(x4==61 && y4==15)||(x4==62 && y4==15)||(x4==2 && y4==16)||(x4==3 && y4==16)||(x4==6 && y4==16)||(x4==7 && y4==16)||(x4==12 && y4==16)||(x4==13 && y4==16)||(x4==14 && y4==16)||(x4==15 && y4==16)||(x4==16 && y4==16)||(x4==17 && y4==16)||(x4==18 && y4==16)||(x4==19 && y4==16)||(x4==20 && y4==16)||(x4==21 && y4==16)||(x4==22 && y4==16)||(x4==23 && y4==16)||(x4==24 && y4==16)||(x4==25 && y4==16)||(x4==26 && y4==16)||(x4==27 && y4==16)||(x4==28 && y4==16)||(x4==29 && y4==16)||(x4==33 && y4==16)||(x4==34 && y4==16)||(x4==35 && y4==16)||(x4==36 && y4==16)||(x4==37 && y4==16)||(x4==38 && y4==16)||(x4==39 && y4==16)||(x4==40 && y4==16)||(x4==41 && y4==16)||(x4==42 && y4==16)||(x4==43 && y4==16)||(x4==44 && y4==16)||(x4==45 && y4==16)||(x4==46 && y4==16)||(x4==47 && y4==16)||(x4==48 && y4==16)||(x4==49 && y4==16)||(x4==50 && y4==16)||(x4==51 && y4==16)||(x4==52 && y4==16)||(x4==53 && y4==16)||(x4==54 && y4==16)||(x4==55 && y4==16)||(x4==56 && y4==16)||(x4==57 && y4==16)||(x4==58 && y4==16)||(x4==59 && y4==16)||(x4==60 && y4==16)||(x4==61 && y4==16)||(x4==62 && y4==16)||(x4==2 && y4==17)||(x4==6 && y4==17)||(x4==7 && y4==17)||(x4==39 && y4==17)||(x4==40 && y4==17)||(x4==41 && y4==17)||(x4==6 && y4==18)||(x4==7 && y4==18)||(x4==39 && y4==18)||(x4==40 && y4==18)||(x4==6 && y4==19)||(x4==7 && y4==19)||(x4==38 && y4==19)||(x4==39 && y4==19)||(x4==40 && y4==19)||(x4==6 && y4==20)||(x4==7 && y4==20)||(x4==12 && y4==20)||(x4==13 && y4==20)||(x4==14 && y4==20)||(x4==15 && y4==20)||(x4==16 && y4==20)||(x4==17 && y4==20)||(x4==18 && y4==20)||(x4==19 && y4==20)||(x4==20 && y4==20)||(x4==21 && y4==20)||(x4==22 && y4==20)||(x4==23 && y4==20)||(x4==24 && y4==20)||(x4==25 && y4==20)||(x4==26 && y4==20)||(x4==27 && y4==20)||(x4==28 && y4==20)||(x4==29 && y4==20)||(x4==38 && y4==20)||(x4==39 && y4==20)||(x4==40 && y4==20)||(x4==41 && y4==20)||(x4==42 && y4==20)||(x4==43 && y4==20)||(x4==44 && y4==20)||(x4==45 && y4==20)||(x4==46 && y4==20)||(x4==47 && y4==20)||(x4==48 && y4==20)||(x4==49 && y4==20)||(x4==50 && y4==20)||(x4==51 && y4==20)||(x4==52 && y4==20)||(x4==53 && y4==20)||(x4==54 && y4==20)||(x4==55 && y4==20)||(x4==56 && y4==20)||(x4==57 && y4==20)||(x4==58 && y4==20)||(x4==6 && y4==21)||(x4==7 && y4==21)||(x4==12 && y4==21)||(x4==13 && y4==21)||(x4==14 && y4==21)||(x4==15 && y4==21)||(x4==16 && y4==21)||(x4==17 && y4==21)||(x4==18 && y4==21)||(x4==19 && y4==21)||(x4==20 && y4==21)||(x4==21 && y4==21)||(x4==22 && y4==21)||(x4==23 && y4==21)||(x4==24 && y4==21)||(x4==25 && y4==21)||(x4==26 && y4==21)||(x4==27 && y4==21)||(x4==28 && y4==21)||(x4==29 && y4==21)||(x4==38 && y4==21)||(x4==39 && y4==21)||(x4==40 && y4==21)||(x4==41 && y4==21)||(x4==42 && y4==21)||(x4==43 && y4==21)||(x4==44 && y4==21)||(x4==45 && y4==21)||(x4==46 && y4==21)||(x4==47 && y4==21)||(x4==48 && y4==21)||(x4==49 && y4==21)||(x4==50 && y4==21)||(x4==51 && y4==21)||(x4==52 && y4==21)||(x4==53 && y4==21)||(x4==54 && y4==21)||(x4==55 && y4==21)||(x4==56 && y4==21)||(x4==57 && y4==21)||(x4==58 && y4==21)||(x4==6 && y4==22)||(x4==7 && y4==22)||(x4==12 && y4==22)||(x4==13 && y4==22)||(x4==14 && y4==22)||(x4==27 && y4==22)||(x4==28 && y4==22)||(x4==29 && y4==22)||(x4==56 && y4==22)||(x4==57 && y4==22)||(x4==58 && y4==22)||(x4==6 && y4==23)||(x4==7 && y4==23)||(x4==12 && y4==23)||(x4==13 && y4==23)||(x4==14 && y4==23)||(x4==27 && y4==23)||(x4==28 && y4==23)||(x4==29 && y4==23)||(x4==56 && y4==23)||(x4==57 && y4==23)||(x4==58 && y4==23)||(x4==6 && y4==24)||(x4==7 && y4==24)||(x4==12 && y4==24)||(x4==13 && y4==24)||(x4==14 && y4==24)||(x4==27 && y4==24)||(x4==28 && y4==24)||(x4==29 && y4==24)||(x4==56 && y4==24)||(x4==57 && y4==24)||(x4==6 && y4==25)||(x4==7 && y4==25)||(x4==12 && y4==25)||(x4==13 && y4==25)||(x4==14 && y4==25)||(x4==27 && y4==25)||(x4==28 && y4==25)||(x4==29 && y4==25)||(x4==56 && y4==25)||(x4==57 && y4==25)||(x4==6 && y4==26)||(x4==7 && y4==26)||(x4==12 && y4==26)||(x4==13 && y4==26)||(x4==14 && y4==26)||(x4==27 && y4==26)||(x4==28 && y4==26)||(x4==29 && y4==26)||(x4==55 && y4==26)||(x4==56 && y4==26)||(x4==57 && y4==26)||(x4==6 && y4==27)||(x4==7 && y4==27)||(x4==12 && y4==27)||(x4==13 && y4==27)||(x4==14 && y4==27)||(x4==15 && y4==27)||(x4==16 && y4==27)||(x4==17 && y4==27)||(x4==18 && y4==27)||(x4==19 && y4==27)||(x4==20 && y4==27)||(x4==21 && y4==27)||(x4==22 && y4==27)||(x4==23 && y4==27)||(x4==24 && y4==27)||(x4==25 && y4==27)||(x4==26 && y4==27)||(x4==27 && y4==27)||(x4==28 && y4==27)||(x4==29 && y4==27)||(x4==54 && y4==27)||(x4==55 && y4==27)||(x4==56 && y4==27)||(x4==57 && y4==27)||(x4==6 && y4==28)||(x4==7 && y4==28)||(x4==12 && y4==28)||(x4==13 && y4==28)||(x4==14 && y4==28)||(x4==15 && y4==28)||(x4==16 && y4==28)||(x4==17 && y4==28)||(x4==18 && y4==28)||(x4==19 && y4==28)||(x4==20 && y4==28)||(x4==21 && y4==28)||(x4==22 && y4==28)||(x4==23 && y4==28)||(x4==24 && y4==28)||(x4==25 && y4==28)||(x4==26 && y4==28)||(x4==27 && y4==28)||(x4==28 && y4==28)||(x4==29 && y4==28)||(x4==45 && y4==28)||(x4==46 && y4==28)||(x4==47 && y4==28)||(x4==48 && y4==28)||(x4==49 && y4==28)||(x4==50 && y4==28)||(x4==51 && y4==28)||(x4==52 && y4==28)||(x4==53 && y4==28)||(x4==54 && y4==28)||(x4==55 && y4==28)||(x4==56 && y4==28)||(x4==6 && y4==29)||(x4==7 && y4==29)||(x4==12 && y4==29)||(x4==13 && y4==29)||(x4==14 && y4==29)||(x4==27 && y4==29)||(x4==28 && y4==29)||(x4==29 && y4==29)||(x4==45 && y4==29)||(x4==46 && y4==29)||(x4==47 && y4==29)||(x4==48 && y4==29)||(x4==49 && y4==29)||(x4==50 && y4==29)||(x4==51 && y4==29)||(x4==52 && y4==29)||(x4==53 && y4==29)||(x4==54 && y4==29)||(x4==55 && y4==29)||(x4==5 && y4==30)||(x4==6 && y4==30)||(x4==7 && y4==30)||(x4==12 && y4==30)||(x4==13 && y4==30)||(x4==14 && y4==30)||(x4==27 && y4==30)||(x4==28 && y4==30)||(x4==29 && y4==30)))	
				// Width: 64, Height: 32 From: /home/wanncy/����/image2verilog/signal.png
			begin {red,green,blue} <= 12'b1111_1111_1111; end
			else begin {red,green,blue} <= 12'b0000_0000_0000; end			
			end
			
			end
		else if(game_status == `Over)
			begin
			x <= (x_pix - 300 + 50);
			y <= (y_pix - 200 + 8);
			if((x==3 && y==1)||(x==4 && y==1)||(x==5 && y==1)||(x==9 && y==1)||(x==10 && y==1)||(x==11 && y==1)||(x==59 && y==1)||(x==60 && y==1)||(x==61 && y==1)||(x==65 && y==1)||(x==66 && y==1)||(x==2 && y==2)||(x==3 && y==2)||(x==58 && y==2)||(x==59 && y==2)||(x==66 && y==2)||(x==67 && y==2)||(x==1 && y==3)||(x==2 && y==3)||(x==57 && y==3)||(x==58 && y==3)||(x==66 && y==3)||(x==67 && y==3)||(x==1 && y==4)||(x==2 && y==4)||(x==16 && y==4)||(x==17 && y==4)||(x==18 && y==4)||(x==19 && y==4)||(x==20 && y==4)||(x==24 && y==4)||(x==25 && y==4)||(x==26 && y==4)||(x==27 && y==4)||(x==29 && y==4)||(x==30 && y==4)||(x==31 && y==4)||(x==32 && y==4)||(x==34 && y==4)||(x==35 && y==4)||(x==36 && y==4)||(x==37 && y==4)||(x==44 && y==4)||(x==45 && y==4)||(x==46 && y==4)||(x==47 && y==4)||(x==48 && y==4)||(x==57 && y==4)||(x==58 && y==4)||(x==66 && y==4)||(x==67 && y==4)||(x==69 && y==4)||(x==70 && y==4)||(x==71 && y==4)||(x==72 && y==4)||(x==78 && y==4)||(x==79 && y==4)||(x==84 && y==4)||(x==85 && y==4)||(x==86 && y==4)||(x==87 && y==4)||(x==88 && y==4)||(x==90 && y==4)||(x==91 && y==4)||(x==92 && y==4)||(x==93 && y==4)||(x==96 && y==4)||(x==97 && y==4)||(x==98 && y==4)||(x==1 && y==5)||(x==14 && y==5)||(x==15 && y==5)||(x==16 && y==5)||(x==19 && y==5)||(x==20 && y==5)||(x==23 && y==5)||(x==24 && y==5)||(x==26 && y==5)||(x==27 && y==5)||(x==28 && y==5)||(x==29 && y==5)||(x==31 && y==5)||(x==32 && y==5)||(x==33 && y==5)||(x==34 && y==5)||(x==36 && y==5)||(x==37 && y==5)||(x==43 && y==5)||(x==44 && y==5)||(x==47 && y==5)||(x==48 && y==5)||(x==56 && y==5)||(x==57 && y==5)||(x==66 && y==5)||(x==67 && y==5)||(x==68 && y==5)||(x==69 && y==5)||(x==71 && y==5)||(x==72 && y==5)||(x==78 && y==5)||(x==79 && y==5)||(x==83 && y==5)||(x==84 && y==5)||(x==87 && y==5)||(x==88 && y==5)||(x==89 && y==5)||(x==90 && y==5)||(x==92 && y==5)||(x==93 && y==5)||(x==94 && y==5)||(x==95 && y==5)||(x==96 && y==5)||(x==1 && y==6)||(x==5 && y==6)||(x==6 && y==6)||(x==7 && y==6)||(x==8 && y==6)||(x==9 && y==6)||(x==10 && y==6)||(x==13 && y==6)||(x==14 && y==6)||(x==19 && y==6)||(x==20 && y==6)||(x==26 && y==6)||(x==27 && y==6)||(x==28 && y==6)||(x==31 && y==6)||(x==32 && y==6)||(x==33 && y==6)||(x==36 && y==6)||(x==37 && y==6)||(x==42 && y==6)||(x==43 && y==6)||(x==47 && y==6)||(x==48 && y==6)||(x==56 && y==6)||(x==57 && y==6)||(x==66 && y==6)||(x==67 && y==6)||(x==71 && y==6)||(x==72 && y==6)||(x==73 && y==6)||(x==77 && y==6)||(x==78 && y==6)||(x==82 && y==6)||(x==83 && y==6)||(x==87 && y==6)||(x==88 && y==6)||(x==92 && y==6)||(x==93 && y==6)||(x==94 && y==6)||(x==1 && y==7)||(x==4 && y==7)||(x==5 && y==7)||(x==8 && y==7)||(x==9 && y==7)||(x==10 && y==7)||(x==13 && y==7)||(x==14 && y==7)||(x==18 && y==7)||(x==19 && y==7)||(x==20 && y==7)||(x==26 && y==7)||(x==27 && y==7)||(x==28 && y==7)||(x==31 && y==7)||(x==32 && y==7)||(x==33 && y==7)||(x==36 && y==7)||(x==37 && y==7)||(x==41 && y==7)||(x==42 && y==7)||(x==45 && y==7)||(x==46 && y==7)||(x==47 && y==7)||(x==56 && y==7)||(x==57 && y==7)||(x==65 && y==7)||(x==66 && y==7)||(x==72 && y==7)||(x==73 && y==7)||(x==76 && y==7)||(x==77 && y==7)||(x==81 && y==7)||(x==82 && y==7)||(x==85 && y==7)||(x==86 && y==7)||(x==87 && y==7)||(x==92 && y==7)||(x==93 && y==7)||(x==94 && y==7)||(x==1 && y==8)||(x==8 && y==8)||(x==9 && y==8)||(x==12 && y==8)||(x==13 && y==8)||(x==17 && y==8)||(x==18 && y==8)||(x==19 && y==8)||(x==25 && y==8)||(x==26 && y==8)||(x==27 && y==8)||(x==31 && y==8)||(x==32 && y==8)||(x==35 && y==8)||(x==36 && y==8)||(x==41 && y==8)||(x==42 && y==8)||(x==43 && y==8)||(x==44 && y==8)||(x==45 && y==8)||(x==56 && y==8)||(x==57 && y==8)||(x==65 && y==8)||(x==66 && y==8)||(x==72 && y==8)||(x==73 && y==8)||(x==75 && y==8)||(x==76 && y==8)||(x==81 && y==8)||(x==82 && y==8)||(x==83 && y==8)||(x==84 && y==8)||(x==85 && y==8)||(x==91 && y==8)||(x==92 && y==8)||(x==93 && y==8)||(x==1 && y==9)||(x==2 && y==9)||(x==7 && y==9)||(x==8 && y==9)||(x==9 && y==9)||(x==12 && y==9)||(x==13 && y==9)||(x==16 && y==9)||(x==17 && y==9)||(x==18 && y==9)||(x==19 && y==9)||(x==25 && y==9)||(x==26 && y==9)||(x==30 && y==9)||(x==31 && y==9)||(x==35 && y==9)||(x==36 && y==9)||(x==41 && y==9)||(x==42 && y==9)||(x==56 && y==9)||(x==57 && y==9)||(x==58 && y==9)||(x==64 && y==9)||(x==65 && y==9)||(x==72 && y==9)||(x==73 && y==9)||(x==74 && y==9)||(x==75 && y==9)||(x==81 && y==9)||(x==82 && y==9)||(x==91 && y==9)||(x==92 && y==9)||(x==1 && y==10)||(x==2 && y==10)||(x==3 && y==10)||(x==7 && y==10)||(x==8 && y==10)||(x==9 && y==10)||(x==12 && y==10)||(x==13 && y==10)||(x==15 && y==10)||(x==16 && y==10)||(x==17 && y==10)||(x==18 && y==10)||(x==19 && y==10)||(x==20 && y==10)||(x==21 && y==10)||(x==22 && y==10)||(x==25 && y==10)||(x==26 && y==10)||(x==30 && y==10)||(x==31 && y==10)||(x==35 && y==10)||(x==36 && y==10)||(x==38 && y==10)||(x==39 && y==10)||(x==41 && y==10)||(x==42 && y==10)||(x==47 && y==10)||(x==48 && y==10)||(x==57 && y==10)||(x==58 && y==10)||(x==62 && y==10)||(x==63 && y==10)||(x==64 && y==10)||(x==72 && y==10)||(x==73 && y==10)||(x==74 && y==10)||(x==81 && y==10)||(x==82 && y==10)||(x==87 && y==10)||(x==88 && y==10)||(x==91 && y==10)||(x==92 && y==10)||(x==2 && y==11)||(x==3 && y==11)||(x==4 && y==11)||(x==5 && y==11)||(x==6 && y==11)||(x==7 && y==11)||(x==8 && y==11)||(x==9 && y==11)||(x==12 && y==11)||(x==13 && y==11)||(x==14 && y==11)||(x==15 && y==11)||(x==18 && y==11)||(x==19 && y==11)||(x==20 && y==11)||(x==24 && y==11)||(x==25 && y==11)||(x==26 && y==11)||(x==30 && y==11)||(x==31 && y==11)||(x==35 && y==11)||(x==36 && y==11)||(x==37 && y==11)||(x==38 && y==11)||(x==42 && y==11)||(x==43 && y==11)||(x==44 && y==11)||(x==45 && y==11)||(x==46 && y==11)||(x==47 && y==11)||(x==58 && y==11)||(x==59 && y==11)||(x==60 && y==11)||(x==61 && y==11)||(x==62 && y==11)||(x==63 && y==11)||(x==72 && y==11)||(x==73 && y==11)||(x==82 && y==11)||(x==83 && y==11)||(x==84 && y==11)||(x==85 && y==11)||(x==86 && y==11)||(x==87 && y==11)||(x==91 && y==11)||(x==92 && y==11)||(x==7 && y==12)||(x==8 && y==12)||(x==1 && y==13)||(x==2 && y==13)||(x==6 && y==13)||(x==7 && y==13)||(x==1 && y==14)||(x==2 && y==14)||(x==3 && y==14)||(x==4 && y==14)||(x==5 && y==14)||(x==6 && y==14)) begin {red,green,blue} <= 12'b1111_1111_1111; end
			else begin {red,green,blue} <= 12'b0000_0000_0000; end// Width: 99, Height: 15 From: /home/wanncy/图片/game_over.png	
			end
	end
		
endmodule

